/*
 * File based on : MParygin/v.vga.font8x16 (Github)
 * 
 * This file implements a Character ROM for translating ASCII
 * character codes into 8x16 pixel image.
 *
 * The input to the module is:
 *  1) 8 bit ASCII code,
 *  2) column select, 0..7, which indicates which of the 8 pixels of the character
 *     image will be returned
 *  3) row select, 0..15, which indicates which of the 16 rows of pixels of the character
 *     image will be returned
 */

module AnalyzerFont (
	input	clk,
	input	[2:0]	col,
	input	[3:0]	row,
	input	[7:0]	ascii,
	output	pixel
);

reg[128:0] char;
wire[7:0] pix_addr;
		 
always@(clk)
begin
	case (ascii)
      8'h00 : char = 128'h00000000000000000000000000000000;
		8'h01 : char = 128'h000000007e818199bd8181a5817e0000;
	   8'h02 : char = 128'h000000007effffe7c3ffffdbff7e0000;
		8'h03 : char = 128'h0000000010387cfefefefe6c00000000;
		8'h04 : char = 128'h000000000010387cfe7c381000000000;
		8'h05 : char = 128'h000000003c1818e7e7e73c3c18000000;
		8'h06 : char = 128'h000000003c18187effff7e3c18000000;
		8'h07 : char = 128'h000000003c1818e7e7e73c3c18000000;
		8'h08 : char = 128'hffffffffffffe7c3c3e7ffffffffffff;
		8'h09 : char = 128'h00000000003c664242663c0000000000;
		8'h0A : char = 128'hffffffffffc399bdbd99c3ffffffffff;
		8'h0B : char = 128'h0000000078cccccccc78321a0e1e0000;
		8'h0C : char = 128'h0000000018187e183c666666663c0000;
		8'h0D : char = 128'h00000000e0f070303030303f333f0000;
		8'h0E : char = 128'h000000c0e6e767636363637f637f0000;
		8'h0F : char = 128'h000000001818db3ce73cdb1818000000;
		
		8'h10 : char = 128'h0000000080c0e0f0f8fef8f0e0c08000;
		8'h11 : char = 128'h0000000002060e1e3efe3e1e0e060200;
		8'h12 : char = 128'h0000000000183c7e1818187e3c180000;
		8'h13 : char = 128'h00000000666600666666666666660000;
		8'h14 : char = 128'h000000001b1b1b1b1b7bdbdbdb7f0000;
		8'h15 : char = 128'h0000007cc60c386cc6c66c3860c67c00;
		8'h16 : char = 128'h00000000fefefefe0000000000000000;
	   8'h17 : char = 128'h000000007e183c7e1818187e3c180000;
		8'h18 : char = 128'h00000000181818181818187e3c180000;
		8'h19 : char = 128'h00000000183c7e181818181818180000;
		8'h1A : char = 128'h000000000000180cfe0c180000000000;
		8'h1B : char = 128'h0000000000003060fe60300000000000;
		8'h1C : char = 128'h000000000000fec0c0c0000000000000;
		8'h1D : char = 128'h0000000000002466ff66240000000000;
		8'h1E : char = 128'h0000000000fefe7c7c38381000000000;
		8'h1F : char = 128'h00000000001038387c7cfefe00000000;
				
		8'h20 : char = 128'h00000000000000000000000000000000;
		8'h21 : char = 128'h000000001818001818183c3c3c180000;
		8'h22 : char = 128'h00000000000000000000002466666600;
		8'h23 : char = 128'h000000006c6cfe6c6c6cfe6c6c000000;
		8'h24 : char = 128'h000018187cc68606067cc0c2c67c1818;
		8'h25 : char = 128'h0000000086c66030180cc6c200000000;
		8'h26 : char = 128'h0000000076ccccccdc76386c6c380000;
		8'h27 : char = 128'h00000000000000000000006030303000;
		8'h28 : char = 128'h000000000c18303030303030180c0000;
		8'h29 : char = 128'h0000000030180c0c0c0c0c0c18300000;
		8'h2A : char = 128'h000000000000663cff3c660000000000;
		8'h2B : char = 128'h00000000000018187e18180000000000;
		8'h2C : char = 128'h00000030181818000000000000000000;
		8'h2D : char = 128'h00000000000000007e00000000000000;
		8'h2E : char = 128'h00000000181800000000000000000000;
		8'h2F : char = 128'h0000000080c06030180c060200000000;
		
		8'h30 : char = 128'h000000007cc6c6e6f6decec6c67c0000;
		8'h31 : char = 128'h000000007e1818181818187838180000;
		8'h32 : char = 128'h00000000fec6c06030180c06c67c0000;
		8'h33 : char = 128'h000000007cc60606063c0606c67c0000;
		8'h34 : char = 128'h000000001e0c0c0cfecc6c3c1c0c0000;
		8'h35 : char = 128'h000000007cc6060606fcc0c0c0fe0000;
		8'h36 : char = 128'h000000007cc6c6c6c6fcc0c060380000;
		8'h37 : char = 128'h0000000030303030180c0606c6fe0000;
		8'h38 : char = 128'h000000007cc6c6c6c67cc6c6c67c0000;
		8'h39 : char = 128'h00000000780c0606067ec6c6c67c0000;
		8'h3A : char = 128'h00000000001818000000181800000000;
		8'h3B : char = 128'h00000000301818000000181800000000;
		8'h3C : char = 128'h00000000060c18306030180c06000000;
		8'h3D : char = 128'h000000000000007e00007e0000000000;
		8'h3E : char = 128'h000000006030180c060c183060000000;
		8'h3F : char = 128'h000000001818001818180cc6c67c0000;
			
		8'h40 : char = 128'h000000007cc0dcdededec6c6c67c0000;
		8'h41 : char = 128'h00000000c6c6c6c6fec6c66c38100000;
		8'h42 : char = 128'h00000000fc666666667c666666fc0000;
		8'h43 : char = 128'h000000003c66c2c0c0c0c0c2663c0000;
		8'h44 : char = 128'h00000000f86c6666666666666cf80000;
		8'h45 : char = 128'h00000000fe6662606878686266fe0000;
		8'h46 : char = 128'h00000000f06060606878686266fe0000;
		8'h47 : char = 128'h000000003a66c6c6dec0c0c2663c0000;
		8'h48 : char = 128'h00000000c6c6c6c6c6fec6c6c6c60000;
		8'h49 : char = 128'h000000003c18181818181818183c0000;
		8'h4A : char = 128'h0000000078cccccc0c0c0c0c0c1e0000;
		8'h4B : char = 128'h00000000e666666c78786c6666e60000;
		8'h4C : char = 128'h00000000fe6662606060606060f00000;
		8'h4D : char = 128'h00000000c3c3c3c3c3dbffffe7c30000;
		8'h4E : char = 128'h00000000c6c6c6c6cedefef6e6c60000;
		8'h4F : char = 128'h000000007cc6c6c6c6c6c6c6c67c0000;
		
		8'h50 : char = 128'h00000000f0606060607c666666fc0000;
		8'h51 : char = 128'h00000e0c7cded6c6c6c6c6c6c67c0000;
		8'h52 : char = 128'h00000000e66666666c7c666666fc0000;
		8'h53 : char = 128'h000000007cc6c6060c3860c6c67c0000;
		8'h54 : char = 128'h000000003c18181818181899dbff0000;
		8'h55 : char = 128'h000000007cc6c6c6c6c6c6c6c6c60000;
		8'h56 : char = 128'h00000000183c66c3c3c3c3c3c3c30000;
		8'h57 : char = 128'h000000006666ffdbdbc3c3c3c3c30000;
		8'h58 : char = 128'h00000000c3c3663c18183c66c3c30000;
		8'h59 : char = 128'h000000003c181818183c66c3c3c30000;
		8'h5A : char = 128'h00000000ffc3c16030180c86c3ff0000;
		8'h5B : char = 128'h000000003c30303030303030303c0000;
		8'h5C : char = 128'h0000000002060e1c3870e0c080000000;
		8'h5D : char = 128'h000000003c0c0c0c0c0c0c0c0c3c0000;
		8'h5E : char = 128'h000000000000000000000000c66c3810;
		8'h5F : char = 128'h0000ff00000000000000000000000000;
				
		8'h60 : char = 128'h00000000000000000000000000183030;
		8'h61 : char = 128'h0000000076cccccc7c0c780000000000;
		8'h62 : char = 128'h000000007c666666666c786060e00000;
		8'h63 : char = 128'h000000007cc6c0c0c0c67c0000000000;
		8'h64 : char = 128'h0000000076cccccccc6c3c0c0c1c0000;
		8'h65 : char = 128'h000000007cc6c0c0fec67c0000000000;
		8'h66 : char = 128'h00000000f060606060f060646c380000;
		8'h67 : char = 128'h0078cc0c7ccccccccccc760000000000;
		8'h68 : char = 128'h00000000e666666666766c6060e00000;
		8'h69 : char = 128'h000000003c1818181818380018180000;
		8'h6A : char = 128'h003c66660606060606060e0006060000;
		8'h6B : char = 128'h00000000e6666c78786c666060e00000;
		8'h6C : char = 128'h000000003c1818181818181818380000;
		8'h6D : char = 128'h00000000dbdbdbdbdbffe60000000000;
		8'h6E : char = 128'h00000000666666666666dc0000000000;
		8'h6F : char = 128'h000000007cc6c6c6c6c67c0000000000;
		
		8'h70 : char = 128'h00f060607c6666666666dc0000000000;
		8'h71 : char = 128'h001e0c0c7ccccccccccc760000000000;
		8'h72 : char = 128'h00000000f06060606676dc0000000000;
		8'h73 : char = 128'h000000007cc60c3860c67c0000000000;
		8'h74 : char = 128'h000000001c3630303030fc3030100000;
		8'h75 : char = 128'h0000000076cccccccccccc0000000000;
		8'h76 : char = 128'h00000000183c66c3c3c3c30000000000;
		8'h77 : char = 128'h0000000066ffdbdbc3c3c30000000000;
		8'h78 : char = 128'h00000000c3663c183c66c30000000000;
		8'h79 : char = 128'h00f80c067ec6c6c6c6c6c60000000000;
		8'h7A : char = 128'h00000000fec6603018ccfe0000000000;
		8'h7B : char = 128'h000000000e18181818701818180e0000;
		8'h7C : char = 128'h00000000181818181800181818180000;
		8'h7D : char = 128'h0000000070181818180e181818700000;
		8'h7E : char = 128'h000000000000000000000000dc760000;
		8'h7F : char = 128'h0000000000fec6c6c66c381000000000;
				
		8'h80 : char = 128'h00007c060c3c66c2c0c0c0c2663c0000;
		8'h81 : char = 128'h0000000076cccccccccccc0000cc0000;
		8'h82 : char = 128'h000000007cc6c0c0fec67c0030180c00;
		8'h83 : char = 128'h0000000076cccccc7c0c78006c381000;
		8'h84 : char = 128'h0000000076cccccc7c0c780000cc0000;
		8'h85 : char = 128'h0000000076cccccc7c0c780018306000;
		8'h86 : char = 128'h0000000076cccccc7c0c7800386c3800;
		8'h87 : char = 128'h0000003c060c3c666060663c00000000;
		8'h88 : char = 128'h000000007cc6c0c0fec67c006c381000;
		8'h89 : char = 128'h000000007cc6c0c0fec67c0000c60000;
		8'h8A : char = 128'h000000007cc6c0c0fec67c0018306000;
		8'h8B : char = 128'h000000003c1818181818380000660000;
		8'h8C : char = 128'h000000003c18181818183800663c1800;
		8'h8D : char = 128'h000000003c1818181818380018306000;
		8'h8E : char = 128'h00000000c6c6c6fec6c66c381000c600;
		8'h8F : char = 128'h00000000c6c6c6fec6c66c3800386c38;
		
		8'h90 : char = 128'h00000000fe6660607c6066fe00603018;
		8'h91 : char = 128'h0000000077dcd87e1b3b6e0000000000;
		8'h92 : char = 128'h00000000ceccccccccfecccc6c3e0000;
		8'h93 : char = 128'h000000007cc6c6c6c6c67c006c381000;
		8'h94 : char = 128'h000000007cc6c6c6c6c67c0000c60000;
		8'h95 : char = 128'h000000007cc6c6c6c6c67c0018306000;
		8'h96 : char = 128'h0000000076cccccccccccc00cc783000;
		8'h97 : char = 128'h0000000076cccccccccccc0018306000;
		8'h98 : char = 128'h00780c067ec6c6c6c6c6c60000c60000;
		8'h99 : char = 128'h000000007cc6c6c6c6c6c6c67c00c600;
		8'h9A : char = 128'h000000007cc6c6c6c6c6c6c6c600c600;
		8'h9B : char = 128'h0000000018187ec3c0c0c0c37e181800;
		8'h9C : char = 128'h00000000fce660606060f060646c3800;
		8'h9D : char = 128'h00000000181818ff18ff183c66c30000;
		8'h9E : char = 128'h00000000f36666666f66627c6666fc00;
		8'h9F : char = 128'h000070d818181818187e1818181b0e00;
				
		8'hA0 : char = 128'h0000000076cccccc7c0c780060301800;
		8'hA1 : char = 128'h000000003c1818181818380030180c00;
		8'hA2 : char = 128'h000000007cc6c6c6c6c67c0060301800;
		8'hA3 : char = 128'h0000000076cccccccccccc0060301800;
		8'hA4 : char = 128'h00000000666666666666dc00dc760000;
		8'hA5 : char = 128'h00000000c6c6c6cedefef6e6c600dc76;
		8'hA6 : char = 128'h0000000000000000007e003e6c6c3c00;
		8'hA7 : char = 128'h0000000000000000007c00386c6c3800;
		8'hA8 : char = 128'h000000007cc6c6c06030300030300000;
		8'hA9 : char = 128'h0000000000c0c0c0c0fe000000000000;
		8'hAA : char = 128'h000000000006060606fe000000000000;
		8'hAB : char = 128'h00001f0c069bce603018ccc6c2c0c000;
		8'hAC : char = 128'h000006063e96ce663018ccc6c2c0c000;
		8'hAD : char = 128'h00000000183c3c3c1818180018180000;
		8'hAE : char = 128'h000000000000366cd86c360000000000;
		8'hAF : char = 128'h000000000000d86c366cd80000000000;
		
		8'hB0 : char = 128'h44114411441144114411441144114411;
		8'hB1 : char = 128'haa55aa55aa55aa55aa55aa55aa55aa55;
		8'hB2 : char = 128'h77dd77dd77dd77dd77dd77dd77dd77dd;
		8'hB3 : char = 128'h18181818181818181818181818181818;
		8'hB4 : char = 128'h1818181818181818f818181818181818;
		8'hB5 : char = 128'h1818181818181818f818f81818181818;
		8'hB6 : char = 128'h3636363636363636f636363636363636;
		8'hB7 : char = 128'h3636363636363636fe00000000000000;
		8'hB8 : char = 128'h1818181818181818f818f80000000000;
		8'hB9 : char = 128'h3636363636363636f606f63636363636;
		8'hBA : char = 128'h36363636363636363636363636363636;
		8'hBB : char = 128'h3636363636363636f606fe0000000000;
		8'hBC : char = 128'h0000000000000000fe06f63636363636;
		8'hBD : char = 128'h0000000000000000fe36363636363636;
		8'hBE : char = 128'h0000000000000000f818f81818181818;
		8'hBF : char = 128'h1818181818181818f800000000000000;
				
		8'hC0 : char = 128'h00000000000000001f18181818181818;
		8'hC1 : char = 128'h0000000000000000ff18181818181818;
		8'hC2 : char = 128'h1818181818181818ff00000000000000;
		8'hC3 : char = 128'h18181818181818181f18181818181818;
		8'hC4 : char = 128'h0000000000000000ff00000000000000;
		8'hC5 : char = 128'h1818181818181818ff18181818181818;
		8'hC6 : char = 128'h18181818181818181f181f1818181818;
		8'hC7 : char = 128'h36363636363636363736363636363636;
		8'hC8 : char = 128'h00000000000000003f30373636363636;
		8'hC9 : char = 128'h363636363636363637303f0000000000;
		8'hCA : char = 128'h0000000000000000ff00f73636363636;
		8'hCB : char = 128'h3636363636363636f700ff0000000000;
		8'hCC : char = 128'h36363636363636363730373636363636;
		8'hCD : char = 128'h0000000000000000ff00ff0000000000;
		8'hCE : char = 128'h3636363636363636f700f73636363636;
		8'hCF : char = 128'h0000000000000000ff00ff1818181818;
		
		8'hD0 : char = 128'h0000000000000000ff36363636363636;
		8'hD1 : char = 128'h1818181818181818ff00ff0000000000;
		8'hD2 : char = 128'h3636363636363636ff00000000000000;
		8'hD3 : char = 128'h00000000000000003f36363636363636;
		8'hD4 : char = 128'h00000000000000001f181f1818181818;
		8'hD5 : char = 128'h18181818181818181f181f0000000000;
		8'hD6 : char = 128'h36363636363636363f00000000000000;
		8'hD7 : char = 128'h3636363636363636ff36363636363636;
		8'hD8 : char = 128'h1818181818181818ff18ff1818181818;
		8'hD9 : char = 128'h0000000000000000f818181818181818;
		8'hDA : char = 128'h18181818181818181f00000000000000;
		8'hDB : char = 128'hffffffffffffffffffffffffffffffff;
		8'hDC : char = 128'hffffffffffffffffff00000000000000;
		8'hDD : char = 128'hf0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0;
		8'hDE : char = 128'h0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f;
		8'hDF : char = 128'h000000000000000000ffffffffffffff;
				
		8'hE0 : char = 128'h0000000076dcd8d8d8dc760000000000;
		8'hE1 : char = 128'h00000000ccc6c6c6ccd8cccccc780000;
		8'hE2 : char = 128'h00000000c0c0c0c0c0c0c0c6c6fe0000;
		8'hE3 : char = 128'h000000006c6c6c6c6c6c6cfe00000000;
		8'hE4 : char = 128'h00000000fec66030183060c6fe000000;
		8'hE5 : char = 128'h0000000070d8d8d8d8d87e0000000000;
		8'hE6 : char = 128'h000000c060607c666666666600000000;
		8'hE7 : char = 128'h00000000181818181818dc7600000000;
		8'hE8 : char = 128'h000000007e183c6666663c187e000000;
		8'hE9 : char = 128'h00000000386cc6c6fec6c66c38000000;
		8'hEA : char = 128'h00000000ee6c6c6c6cc6c6c66c380000;
		8'hEB : char = 128'h000000003c666666663e0c18301e0000;
		8'hEC : char = 128'h0000000000007edbdbdb7e0000000000;
		8'hED : char = 128'h00000000c0607ef3dbdb7e0603000000;
		8'hEE : char = 128'h000000001c306060607c6060301c0000;
		8'hEF : char = 128'h00000000c6c6c6c6c6c6c6c67c000000;
		
		8'hF0 : char = 128'h0000000000fe0000fe0000fe00000000;
		8'hF1 : char = 128'h00000000ff000018187e181800000000;
		8'hF2 : char = 128'h000000007e0030180c060c1830000000;
		8'hF3 : char = 128'h000000007e000c18306030180c000000;
		8'hF4 : char = 128'h181818181818181818181b1b1b0e0000;
		8'hF5 : char = 128'h0000000070d8d8d81818181818181818;
		8'hF6 : char = 128'h00000000001818007e00181800000000;
		8'hF7 : char = 128'h000000000000dc7600dc760000000000;
		8'hF8 : char = 128'h0000000000000000000000386c6c3800;
		8'hF9 : char = 128'h00000000000000181800000000000000;
		8'hFA : char = 128'h00000000000000180000000000000000;
		8'hFB : char = 128'h000000001c3c6c6cec0c0c0c0c0c0f00;
		8'hFC : char = 128'h0000000000000000006c6c6c6c6cd800;
		8'hFD : char = 128'h000000000000000000f8c86030d87000;
		8'hFE : char = 128'h00000000007c7c7c7c7c7c7c00000000;
		8'hFF : char = 128'h00000000000000000000000000000000;
   endcase
end

assign pix_addr = {row, col};
assign pixel = char[pix_addr];

endmodule 
