-- -----------------------------------------------------------------------
--
-- Syntiac's generic VHDL support files.
--
-- -----------------------------------------------------------------------
-- Copyright 2005-2008 by Peter Wendrich (pwsoft@syntiac.com)
-- http://www.syntiac.com/fpga64.html
--
-- Modified April 2016 by Dar (darfpga@aol.fr) 
-- http://darfpga.blogspot.fr
--   Remove address register when writing
--
-- Modifies Octiber 2017 by Dar 
--   Add init data with defender cmos value
-- -----------------------------------------------------------------------
--
-- gen_rwram.vhd init with Qix cmos value
--
-- -----------------------------------------------------------------------
--
-- generic ram.
--
-- -----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- -----------------------------------------------------------------------

entity qix_cmos_ram is
	generic (
		dWidth : integer :=  8; -- must be  8 for qix_cmos_ram
		aWidth : integer := 10  -- must be 10 for qix_cmos_ram
	);
	port (
		clk  : in std_logic;
		we   : in std_logic;
		addr : in std_logic_vector((aWidth-1) downto 0);
		d    : in std_logic_vector((dWidth-1) downto 0);
		q    : out std_logic_vector((dWidth-1) downto 0)
	);
end entity;

-- -----------------------------------------------------------------------
--    QIX NONVOLATILE CMOS MEMORY MAP (CPU #2 -- Video) $8400-$87ff
--        $86A9 - $86AA:  When CMOS is valid, these bytes are $55AA
--        $86AC - $86C3:  AUDIT TOTALS -- 4 4-bit BCD digits per setting
--                        (All totals default to: 0000)
--                        $86AC: TOTAL PAID CREDITS
--                        $86AE: LEFT COINS
--                        $86B0: CENTER COINS
--                        $86B2: RIGHT COINS
--                        $86B4: PAID CREDITS
--                        $86B6: AWARDED CREDITS
--                        $86B8: % FREE PLAYS
--                        $86BA: MINUTES PLAYED
--                        $86BC: MINUTES AWARDED
--                        $86BE: % FREE TIME
--                        $86C0: AVG. GAME [SEC]
--                        $86C2: HIGH SCORES
--        $86C4 - $86FF:  High scores -- 10 scores/names, consecutive in memory
--                        Six 4-bit BCD digits followed by 3 ascii bytes
--                        (Default: 030000 QIX)
--        $8700        :  LANGUAGE SELECT (Default: $32)
--                        ENGLISH = $32  FRANCAIS = $33  ESPANOL = $34  DEUTSCH = $35
--        $87D9 - $87DF:  COIN SLOT PROGRAMMING -- 2 4-bit BCD digits per setting
--                        $87D9: STANDARD COINAGE SETTING  (Default: 01)
--                        $87DA: COIN MULTIPLIERS LEFT (Default: 01)
--                        $87DB: COIN MULTIPLIERS CENTER (Default: 04)
--                        $87DC: COIN MULTIPLIERS RIGHT (Default: 01)
--                        $87DD: COIN UNITS FOR CREDIT (Default: 01)
--                        $87DE: COIN UNITS FOR BONUS (Default: 00)
--                        $87DF: MINIMUM COINS (Default: 00)
--        $87E0 - $87EA:  LOCATION PROGRAMMING -- 2 4-bit BCD digits per setting
--                        $87E0: BACKUP HSTD [0000] (Default: 03)
--                        $87E1: MAXIMUM CREDITS (Default: 10)
--                        $87E2: NUMBER OF TURNS (Default: 03)
--                        $87E3: THRESHOLD (Default: 75)
--                        $87E4: TIME LINE (Default: 37)
--                        $87E5: DIFFICULTY 1 (Default: 01)
--                        $87E6: DIFFICULTY 2 (Default: 01)
--                        $87E7: DIFFICULTY 3 (Default: 01)
--                        $87E8: DIFFICULTY 4 (Default: 01)
--                        $87E9: ATTRACT SOUND (Default: 01)
--                        $87EA: TABLE MODE (Default: 00)


architecture rtl of qix_cmos_ram is
	subtype addressRange is integer range 0 to ((2**aWidth)-1);
	type ramDef is array(addressRange) of std_logic_vector((dWidth-1) downto 0);
	
	signal ram: ramDef := (
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0000
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0010
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0020
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0030
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0040
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0050
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0060
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0070
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0080
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0090
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00A0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00B0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00C0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00D0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00E0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x00F0
		
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0100
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0110
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0120
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0130
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0140
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0150
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0160
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0170
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0180
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0190
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01A0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01B0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01C0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01D0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01E0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x01F0
		
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0200
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0210
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0220
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0230
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0240
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0250
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0260
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0270
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0280
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0290
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"55", X"AA", X"00", X"00", X"00", X"00", X"00", -- x02A0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x02B0
		X"00", X"00", X"00", X"00", X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", -- x02C0
		X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", -- x02D0
		X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", -- x02E0
		X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", X"03", X"00", X"00", X"51", X"49", X"58", -- x02F0
		
		X"32", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0300
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0310
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0320
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0330
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0340
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0350
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0360
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0370
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0380
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x0390
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x03A0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x03B0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", -- x03C0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"01", X"01", X"04", X"01", X"01", X"00", X"00", -- x03D0
		X"03", X"10", X"03", X"75", X"37", X"01", X"01", X"01", X"01", X"01", X"00", X"00", X"00", X"00", X"00", X"00", -- x03E0
		X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"  -- x03F0

		);
	
	signal rAddrReg : std_logic_vector((aWidth-1) downto 0);
	signal qReg : std_logic_vector((dWidth-1) downto 0);
begin

-- -----------------------------------------------------------------------
-- Memory write
-- -----------------------------------------------------------------------
	process(clk)
	begin
		if rising_edge(clk) then
			if we = '1' then
				ram(to_integer(unsigned(addr))) <= d;
			end if;
		end if;
	end process;
	
-- -----------------------------------------------------------------------
-- Memory read
-- -----------------------------------------------------------------------
process(clk)
	begin
		if rising_edge(clk) then
			q <= ram(to_integer(unsigned(addr)));
		end if;
	end process;
end architecture;

